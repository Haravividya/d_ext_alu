package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "./../UVME/sequence/d_ext_alu_tx.sv"
    `include "./../UVME/agent/d_ext_alu_sequencer.sv"
    `include "./../UVME/sequence/d_ext_alu_base_seq.sv"
    `include "./../UVME/sequence/FADD_D_seq.sv"
    `include "./../UVME/sequence/FSUB_D_seq.sv"
    `include "./../UVME/sequence/FMUL_D_seq.sv"
    `include "./../UVME/sequence/FDIV_D_seq.sv"
    `include "./../UVME/sequence/FSQRT_D_seq.sv"
    `include "./../UVME/sequence/FMADD_D_seq.sv"
    `include "./../UVME/sequence/FMSUB_D_seq.sv"
    `include "./../UVME/sequence/FNMADD_D_seq.sv"
    `include "./../UVME/sequence/FNMSUB_D_seq.sv"
    `include "./../UVME/sequence/FSGNJ_D_seq.sv"
    `include "./../UVME/sequence/FSGNJN_D_seq.sv"
    `include "./../UVME/sequence/FSGNJX_D_seq.sv"
    `include "./../UVME/sequence/FMIN_D_seq.sv"
    `include "./../UVME/sequence/FMAX_D_seq.sv"
    `include "./../UVME/sequence/FLT_D_seq.sv"
    `include "./../UVME/sequence/FEQ_D_seq.sv"
    `include "./../UVME/sequence/FLE_D_seq.sv"
    `include "./../UVME/sequence/FCVT_S_D_seq.sv"
    `include "./../UVME/sequence/FCVT_D_S_seq.sv"
    `include "./../UVME/sequence/FCVT_D_W_seq.sv"
    `include "./../UVME/sequence/FCVT_D_WU_seq.sv"
    `include "./../UVME/sequence/FCVT_W_D_seq.sv"
    `include "./../UVME/sequence/FCVT_WU_D_seq.sv"
    `include "./../UVME/sequence/FCVT_D_L_seq.sv"
    `include "./../UVME/sequence/FCVT_D_LU_seq.sv"
    `include "./../UVME/sequence/FMV_X_D_seq.sv"
    `include "./../UVME/sequence/FMV_D_X_seq.sv"
    `include "./../UVME/sequence/FCVT_L_D_seq.sv"
    `include "./../UVME/sequence/FCVT_LU_D_seq.sv"
    `include "./../UVME/sequence/FCLASS_D_seq.sv"
    
    `include "./../UVME/sequence/zero_seq.sv"
    `include "./../UVME/sequence/one_seq.sv"
    `include "./../UVME/sequence/corner_seq.sv"
    `include "./../UVME/sequence/random_seq.sv"
    `include "./../UVME/sequence/random_instruction_data_seq.sv"
    //`include "./../UVME/sequence/fcvt_sd_covrage.sv"

    `include "./../UVME/agent/d_ext_alu_driver.sv"
    `include "./../UVME/agent/d_ext_alu_monitor.sv"
    `include "./../UVME/agent/d_ext_alu_agent.sv" 
    `include "./../UVME/env/d_ext_alu_sbd.sv"
    `include "./../UVME/env/d_ext_alu_cov.sv" 
    `include "./../UVME/env/d_ext_alu_env.sv"
    `include "./../UVME/tests/d_ext_alu_base_test.sv"
    `include "./../UVME/tests/FADD_D_Test.sv"
    `include "./../UVME/tests/FSUB_D_Test.sv"
    `include "./../UVME/tests/FMUL_D_Test.sv"
    `include "./../UVME/tests/FDIV_D_Test.sv"
    `include "./../UVME/tests/FSQRT_D_Test.sv"
    `include "./../UVME/tests/FMADD_D_Test.sv"
    `include "./../UVME/tests/FMSUB_D_Test.sv"
    `include "./../UVME/tests/FNMADD_D_Test.sv"
    `include "./../UVME/tests/FNMSUB_D_Test.sv"
    `include "./../UVME/tests/FSGNJ_D_Test.sv"
    `include "./../UVME/tests/FSGNJN_D_Test.sv"
    `include "./../UVME/tests/FSGNJX_D_Test.sv"
    `include "./../UVME/tests/FMIN_D_Test.sv"
    `include "./../UVME/tests/FMAX_D_Test.sv"
    `include "./../UVME/tests/FEQ_D_Test.sv"
    `include "./../UVME/tests/FLT_D_Test.sv"
    `include "./../UVME/tests/FLE_D_Test.sv"
    `include "./../UVME/tests/FCVT_S_D_Test.sv"
    `include "./../UVME/tests/FCVT_D_S_Test.sv"
    `include "./../UVME/tests/FCVT_D_W_Test.sv"
    `include "./../UVME/tests/FCVT_D_WU_Test.sv"
    `include "./../UVME/tests/FCVT_W_D_Test.sv"
    `include "./../UVME/tests/FCVT_WU_D_Test.sv"
    `include "./../UVME/tests/FCVT_D_L_Test.sv"
    `include "./../UVME/tests/FCVT_D_LU_Test.sv"
    `include "./../UVME/tests/FMV_X_D_Test.sv"
    `include "./../UVME/tests/FMV_D_X_Test.sv"
    `include "./../UVME/tests/FCVT_L_D_Test.sv"
    `include "./../UVME/tests/FCVT_LU_D_Test.sv"
    `include "./../UVME/tests/FCLASS_D_Test.sv"  
    `include "./../UVME/tests/zero_test.sv" 
    `include "./../UVME/tests/one_test.sv" 
    `include "./../UVME/tests/corner_test.sv"
    `include "./../UVME/tests/random_test.sv"
    `include "./../UVME/tests/random_instruction_data_test.sv"
    //`include "./../UVME/tests/fcvt_sd_coverage_test.sv"
endpackage
