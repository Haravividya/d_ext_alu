class FCVT_D_WU_seq extends uvm_sequence#(d_ext_alu_tx);
  //factory registration
  `uvm_object_utils(FCVT_D_WU_seq)
  //creating sequence item handle
   d_ext_alu_tx tx;

   int scenario;
  // event seq_done;

  //constructor
   function new(string name="FCVT_D_WU_seq");
        super.new(name);
   endfunction
  
  //Build phase
  function build_phase(uvm_phase phase);
        tx = d_ext_alu_tx::type_id::create("tx");
  endfunction
  
  //task body
  task body();

 
         if (scenario == 1) 
         begin

                `uvm_info (get_type_name(),"Starting Scenario 1:fixed value test case", UVM_LOW)
                `uvm_do_with(tx, {
                                    tx.alu_op  == 5'b10100;
                                    tx.int_rs1 == 32'hFFFFFFFF;
                                                                       
                            })
                `uvm_info (get_type_name(),$sformatf("int_rs1=%h",tx.int_rs1), UVM_LOW)

                `uvm_info(get_type_name(), "Starting Scenario 1: fixed test case done", UVM_LOW)
         end
         
       if (scenario == 2)
       // repeat(10)
       for(int i=0;i<200;i++)


        begin

                `uvm_info(get_type_name(), "Starting Scenario 2: Random test case started", UVM_LOW)
                `uvm_do_with(tx, {
                                    tx.alu_op == 5'b10100;
                                    tx.int_rs1[63:32] == 32'h0;            // Upper 32 bits are 0
                                    tx.int_rs1[31:0] inside {[0 : 32'hFFFFFFFF],[0:32'h7FFFFFFF]}; // Lower 32 bits - Unsigned range
                            })

                `uvm_info(get_type_name(), "Starting Scenario 2: Random test case done", UVM_LOW)
                
        end
  endtask
endclass  



