class FSGNJX_D_Test extends d_ext_alu_base_test;

  // Factory registration
     `uvm_component_utils(FSGNJX_D_Test)
      FSGNJX_D_seq fsgnjx_seq;


  // Constructor
  function new(string name = "FSGNJX_D_Test", uvm_component parent = null);
      super.new(name, parent);
      fsgnjx_seq = FSGNJX_D_seq::type_id::create("fsgnjx_seq");
  endfunction

  // Build Phase
  function void build_phase(uvm_phase phase);
      super.build_phase(phase);
  endfunction

  // Run Phase
  task run_phase(uvm_phase phase);
      phase.raise_objection(this);
     `uvm_info(get_full_name(), $sformatf("Inside the XOR-based sign injection  test"), UVM_MEDIUM)
    // begin
      //fsgnjx_seq.scenario = 1;
      //fsgnjx_seq.start(env.agent.sequencer);
         // @(fmul_seq.seq_done);
     //end
// #10;
   // repeat(10)begin
      fsgnjx_seq.scenario = 2;
      fsgnjx_seq.start(env.agent.sequencer);
      //  @(fmul_seq.seq_done);
   // end
  
     `uvm_info(get_type_name(),$sformatf("random XOR-based sign injection scenario 2 is completed"),UVM_MEDIUM)
     `uvm_info(get_full_name(), $sformatf("Inside the    XOR-based sign injection test done"), UVM_MEDIUM)
      #200;
      phase.drop_objection(this);
  endtask

endclass

